arvind
kamal
nain
